`include "pattern_detector.v"
`include "pattern_detector_mealy.v"

module pattern_detector_tb;
    
    reg clk_i;
    reg rst_i;
    reg d_i;
    wire pattern_detected_o;
    reg [7:0] count;
    integer i;

    pattern_detector_mealy pd0
        (
            .clk_i(clk_i),
            .rst_i(rst_i),
            .d_i(d_i),
            .pattern_detected_o(pattern_detected_o)
        );
/*        
    pattern_detector pd0
        (
            .clk_i(clk_i),
            .rst_i(rst_i),
            .d_i(d_i),
            .pattern_detected_o(pattern_detected_o)
        );
*/
    always begin
        #5 clk_i = 0;
        #5 clk_i = 1;
    end

    initial begin
        i = 690*5;
        rst_i = 0;
        count = 0;

        #40; 
        rst_i = 1;
        #1400;
        $finish;
        
    end

    always begin
        #10
        d_i = $random(i);
    end

    always @ (posedge clk_i) begin
        if(rst_i == 0) begin
            count = 0;
        end

        else begin
            if(pattern_detected_o == 1)
                count = count + 1;
        end
    end

    initial begin
        $monitor("d_i=%0d   pattern_detected_o=%0d  count=%0d", d_i, pattern_detected_o, count);
    end

endmodule
